library verilog;
use verilog.vl_types.all;
entity Lab_1_vlg_vec_tst is
end Lab_1_vlg_vec_tst;
