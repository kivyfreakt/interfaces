library verilog;
use verilog.vl_types.all;
entity clk_divider_vlg_vec_tst is
end clk_divider_vlg_vec_tst;
