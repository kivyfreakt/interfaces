library verilog;
use verilog.vl_types.all;
entity spi_vlg_vec_tst is
end spi_vlg_vec_tst;
