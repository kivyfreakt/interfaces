library verilog;
use verilog.vl_types.all;
entity Lab_1_vlg_check_tst is
    port(
        cs              : in     vl_logic;
        mosi            : in     vl_logic;
        sck             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Lab_1_vlg_check_tst;
