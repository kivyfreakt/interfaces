library verilog;
use verilog.vl_types.all;
entity SPImaster_vlg_vec_tst is
end SPImaster_vlg_vec_tst;
